module alu;


endmodule